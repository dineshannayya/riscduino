//////////////////////////////////////////////////////////////////////
////                                                              ////
////  Active low reset synchronization                           ////
////                                                              ////
////  This file is part of the yifive cores project               ////
////  http://www.opencores.org/cores/yifive/                      ////
////                                                              ////
////  Description:                                                ////
////     Synchronize the active low reset to destination clock    ////
////                                                              ////
////  To Do:                                                      ////
////    nothing                                                   ////
////                                                              ////
////  Author(s):                                                  ////
////      - Dinesh Annayya, dinesha@opencores.org                 ////
////                                                              ////
////  Revision :                                                  ////
////     v0:    June 17, 2021, Dinesh A                           ////
////             Initial version                                  ////
////                                                              ////
//////////////////////////////////////////////////////////////////////
////                                                              ////
//// Copyright (C) 2000 Authors and OPENCORES.ORG                 ////
////                                                              ////
//// This source file may be used and distributed without         ////
//// restriction provided that this copyright statement is not    ////
//// removed from the file and that any derivative work contains  ////
//// the original copyright notice and the associated disclaimer. ////
////                                                              ////
//// This source file is free software; you can redistribute it   ////
//// and/or modify it under the terms of the GNU Lesser General   ////
//// Public License as published by the Free Software Foundation; ////
//// either version 2.1 of the License, or (at your option) any   ////
//// later version.                                               ////
////                                                              ////
//// This source is distributed in the hope that it will be       ////
//// useful, but WITHOUT ANY WARRANTY; without even the implied   ////
//// warranty of MERCHANTABILITY or FITNESS FOR A PARTICULAR      ////
//// PURPOSE.  See the GNU Lesser General Public License for more ////
//// details.                                                     ////
////                                                              ////
//// You should have received a copy of the GNU Lesser General    ////
//// Public License along with this source; if not, download it   ////
//// from http://www.opencores.org/lgpl.shtml                     ////
////                                                              ////
//////////////////////////////////////////////////////////////////////

module reset_sync   (
	      scan_mode  ,
              dclk       , // Destination clock domain
	      arst_n     , // active low async reset
              srst_n 
          );

parameter WIDTH = 1;

input    scan_mode  ; // test mode
input    dclk       ; // Destination clock
input    arst_n     ; // Async Reset
input    srst_n     ; // Sync Reset w.r.t dclk


reg      in_data_s  ; // One   Cycle sync 
reg      in_data_2s ; // two   Cycle sync 

assign srst_n =  (scan_mode) ? arst_n : in_data_2s;

always @(negedge arst_n  or posedge dclk)
begin
   if(arst_n == 1'b0)
   begin
      in_data_s  <= 1'b0;
      in_data_2s <= 1'b0;
   end
   else
   begin
      in_data_s  <= 1'b1;
      in_data_2s <= in_data_s;
   end
end


endmodule

module dac_top (Vout0,
    Vout1,
    Vout2,
    Vout3,
    Vref,
    vccd1,
    vssd1,
    DIn0,
    DIn1,
    DIn2,
    DIn3);
 output Vout0;
 output Vout1;
 output Vout2;
 output Vout3;
 input Vref;
 input vccd1;
 input vssd1;
 input [7:0] DIn0;
 input [7:0] DIn1;
 input [7:0] DIn2;
 input [7:0] DIn3;

endmodule
